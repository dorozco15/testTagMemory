library verilog;
use verilog.vl_types.all;
entity TagMemory_vlg_vec_tst is
end TagMemory_vlg_vec_tst;
